**.subckt Ring Oscillator
x1 net2 net4 net1 net3 inv_1
x2 net2 net5 net4 net3 inv_1
x3 net2 net6 net5 net3 inv_1
x4 net2 net7 net6 net3 inv_1
x5 net2 net1 net7 net3 inv_1
**.ends

* expanding   symbol:  /home/harshit/.xschem/inv_1.sym # of pins=4
* sym_path: /home/harshit/.xschem/inv_1.sym
* sch_path: /home/harshit/.xschem/inv_1.sch
.subckt inv_1  Vdd Vout Vin VSS
*.ipin Vdd
*.ipin VSS
*.opin Vout
*.ipin Vin
XM1 Vout Vin VSS VSS sky130_fd_pr__nfet_01v8 L=0.30 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
XM2 Vout Vin Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.30 W=3.0 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=1 m=1
.ends

.end
