**.subckt pmos_char_1v8
XM1 GND net2 net1 net1 sky130_fd_pr__pfet_01v8 L=0.50 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=5 m=5
Vgs net1 net2 1.8
Vds net1 GND 0
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.dc Vds 0 2.2 1m
.save all
.end


**** end user architecture code
**.ends
.GLOBAL GND
.end
