**.subckt untitled-1
**.ends
.end
