**.subckt ringosc_tran
V1 VDD GND 1.8v
x1 VDD vout VSS ringosc
**** begin user architecture code


.lib /usr/local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt



.include /home/harshit/.xschem/ringosc.spice
.tran 1ps 1s uic
.savecurrents
.save all
.end

**** end user architecture code
**.ends
.GLOBAL GND
.end
